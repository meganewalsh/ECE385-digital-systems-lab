/*module title ( input [12:0]  DrawX, DrawY,
			  input Clk,
           output logic  is_title,
			  output logic [1:0] data_R, data_G );

logic [10:0] start_x = 216;
logic [10:0] start_y = 100;
logic [10:0] size_x = 234;
logic [10:0] size_y = 189;

parameter [88451:0] ROM_R = 88452'h4c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c5353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e515353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c515555554f4c4c4c515555554f4c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c525555554e4c4c4c525555554e4c4c4c525555554e4c4c4c535555554e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e524c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c6b868a8a8a88848484868a8a8a88848484868a8a8a88848484868a8a8a8884848487575555514c4c4c5055555c87848484878a8a8a87847b4e51555555504c4c4c515c8a8a87848484878a8a8a87848484878a8a8a87848484878a8a8a87848484878a8a8a87848484878a8a8a8684584c525555554f4c4c4c52628a8a86848484878a8a8a86848484878a8a8a86848484888a8a8a86848484888a7b554f4c4c4c525555554f4e7e84888a8a8a86848484888a8a8a86848484888a8a8a86848484888a8a8a86848484888a8a8a86848484888a75554e4c4c4c535555554e4c4c4c534c4f555555514c4c99fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7615555514c4c4c50555568f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff834c51555555504c4c4c5172ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c5353504e4e4e5153539dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff65b4e4e51535353504e4e62f1ffffffffffffffffffef5f504e4e4e515353535063f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff88534f4e4e4e525353534f6dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffda52525353534f4e4e4e5258d5ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc54e525353534f4e4e4e525353534f55524c4c4c5055559efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6594c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6594c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6594c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8955504c4c4c515555554f6bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffda51525555554f4c4c4c5259d5ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc54c525555554e4c4c4c535555554e4d50545454504d4d9afffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7605454504d4d4d51545467f1ffffffffffffffffffee5a51545454504d4d4d5168f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff834d515454544f4d4d4d5271ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdb584f4d4d4d525454534f52d4ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7534f4d4d4e535454534e4d4d4e534c4f555555514c4c99fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7615555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7615555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7615555514c4c4c50555568f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff834c51555555504c4c4c5172ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c5354514d4d4d5154549dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff65a4d4d51545454504d4d62f1ffffffffffffffffffef60504d4d4d515454545062f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff88544f4d4d4d515454544f6cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffda52525454534f4d4d4e5258d5ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc54e525454534e4d4d4e535454534e55524c4c4c5055559efffffffffffffffffffffefcfdfdfdfdfdfcfcfcfdfdfffffffffffffffffffff6594c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8fffffffffffffffffffffefdfdfdfcfcfcfdfdfdfdfdfcfcfcfdfdfdfdfdfcfcfeffffffffffffffffffff89554f4c4c4c525555554f6bfffffffffffffffffffffffdfdfdfdfcfcfcfdfdfdfdffffffffffffffffffffda50525555554f4c4c4c525ad5fffffffffffffffffffffdfcfcfdfdfdfdfdfcfcfcfdfdfdfdfdfcfcfcfdfdfdffffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffb06b6f7272726f6b6b6b6f81f8fffffffffffffffffff6594c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffffa672726e6b6b6b6f7272726e6b6b6b6f7272726e6b6bceffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdf7572726e6b6b6b70727294ffffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff8e6b6b717272726d6b6b6b717272726d6b6b6b717272e2ffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c5064f1fffffffffffffffffff6594c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbeffffffffffffffffffff8955504c4c4c515555554f6bffffffffffffffffffffdc5955554f4c4c4c5155557affffffffffffffffffffda51525555554f4c4c4c5259d5ffffffffffffffffffff754c4c525555554f4c4c4c525555554e4c4c4c525555ddffffffffffffffffffffc54c525555554e4c4c4c535555554e4d50545454504d4d9affffffffffffffffffffad54504d4d4d51545454505ef1fffffffffffffffffff7605454504d4d4d51545467f1ffffffffffffffffffee5a51545454504d4d4d5168f8ffffffffffffffffffff954d4d51545454504d4d4d51545454504d4d4d515454c0ffffffffffffffffffff834d51545454504d4d4d5171ffffffffffffffffffffdb524d4d515454544f4d4d74ffffffffffffffffffffdb584f4d4d4d525454534f52d4ffffffffffffffffffff7b54534f4d4d4d525454534f4d4d4d525454534f4d4ddbffffffffffffffffffffc7534f4d4d4e535454534e4d4d4e534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555515cf1fffffffffffffffffff7615555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555515cf1fffffffffffffffffff7615555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555515df1fffffffffffffffffff7615555514c4c4c50555568f2ffffffffffffffffffee5950555555504c4c4c5069f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff834c51555555504c4c4c5172ffffffffffffffffffffdb514c4c51555555504c4c73ffffffffffffffffffffdb594f4c4c4c525555554f51d3ffffffffffffffffffff7b55554f4c4c4c525555554f4c4c4c525555554f4c4cdbffffffffffffffffffffc7544f4c4c4c535555544e4c4c4c5354514d4d4d5154549dffffffffffffffffffffa94d51545454504d4d4d5163f1fffffffffffffffffff65a4d4d51545454504d4d62f1ffffffffffffffffffef60504d4d4d515454545062f8ffffffffffffffffffff995454504d4d4d51545454504d4d4d51545454504d4dbeffffffffffffffffffff8854504d4d4d515454544f6cffffffffffffffffffffdc5854544f4d4d4d51545479ffffffffffffffffffffda52525454544f4d4d4d5258d5ffffffffffffffffffff764d4d525454534f4d4d4d525454534f4d4d4d525454ddffffffffffffffffffffc54e525454534e4d4d4e535454534e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c5064f1fffffffffffffffffff6594c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff754c4c535555554e4c4c4c535555554e4c4c4c535555ddffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c5064f1fffffffffffffffffff6594c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff754c4c535555554e4c4c4c535555554e4c4c4c535555ddffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c5064f1fffffffffffffffffff6594c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c505555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbeffffffffffffffffffff8955504c4c4c51555555506bffffffffffffffffffffdc595555504c4c4c5155557affffffffffffffffffffda51525555554f4c4c4c5259d5ffffffffffffffffffff754c4c525555554f4c4c4c525555554f4c4c4c525555ddffffffffffffffffffffc54c525555544e4c4c4c535555544e4d50545454504d4d9affffffffffffffffffffb25d5a5757575b5d5d5d5a66f1fffffffffffffffffff7605454504d4d4d51545467f1ffffffffffffffffffee5a51545454504d4d4d5168f8ffffffffffffffffffff954d4d51545454504d4d4d51545454504d4d4d515454c0ffffffffffffffffffff834d51545454504d4d4d5171ffffffffffffffffffffdb524d4d515454544f4d4d74ffffffffffffffffffffdb584f4d4d4d525454534f52d4ffffffffffffffffffff7b54534f4d4d4d525454534f4d4d4d525454534f4d4ddbffffffffffffffffffffc7534f4d4d4e535454534e4d4d4e534c4f555555514c4c99fffffffffffffffffffff2e2e1e0e0e0e1e2e2e2e1e2fbfffffffffffffffffff7615555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7615555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7615555514c4c4c50555568f2ffffffffffffffffffee5950555555504c4c4c5069f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff834c51555555504c4c4c5172ffffffffffffffffffffdb514c4c51555555504c4c73ffffffffffffffffffffdb594f4c4c4c525555554f51d3ffffffffffffffffffff7b55554f4c4c4c525555554f4c4c4c525555554f4c4cdbffffffffffffffffffffc7544f4c4c4c535555544e4c4c4c5354514d4d4d5054549dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff65a4d4d51545454504d4d62f1ffffffffffffffffffef60504d4d4d515454545062f8ffffffffffffffffffff9a5454504d4d4d51545454504d4d4d51545454504d4dbeffffffffffffffffffff88544f4d4d4d525454544f6cffffffffffffffffffffdc5854544f4d4d4d52545479ffffffffffffffffffffda51525454544f4d4d4d5259d5ffffffffffffffffffff754d4d535454544e4d4d4d535454544e4d4d4d535454ddffffffffffffffffffffc54d535454544e4d4d4d535454544e55524c4c4c5055559efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6594c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff754c4c535555554e4c4c4c535555554e4c4c4c535555ddffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6594c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff754c4c535555554e4c4c4c535555554e4c4c4c535555ddffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6594c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c505555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbeffffffffffffffffffff8955504c4c4c51555555506bffffffffffffffffffffdc595555504c4c4c5155557affffffffffffffffffffda51525555554f4c4c4c5259d5ffffffffffffffffffff754c4c525555554f4c4c4c525555554f4c4c4c525555ddffffffffffffffffffffc54c525555544e4c4c4c535555544e4d50545454514d4d9afffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7615454504d4d4d51545468f1ffffffffffffffffffee5951545454504d4d4d5168f8ffffffffffffffffffff954d4d51545454504d4d4d51545454504d4d4d515454c0ffffffffffffffffffff834d525454544f4d4d4d5272ffffffffffffffffffffdb514d4d525454544f4d4d73ffffffffffffffffffffdb584f4d4d4d525454544f52d4ffffffffffffffffffff7b54544e4d4d4d535454544e4d4d4d535454544e4d4ddbffffffffffffffffffffc7544e4d4d4d535454544e4d4d4d534c4f555555514c4c99fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7615555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7615555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99fffffffffffffffffffffefdfdfcfcfcfdfdfdfdfdfcfcfcfdfdfdfdfdfcfcfcf5615555514c4c4c50555568f2ffffffffffffffffffee5950555555504c4c4c5069f8ffffffffffffffffffff974f4f53575757524f4f4f53575757524f4f4f535757c1ffffffffffffffffffff834c51555555504c4c4c5172ffffffffffffffffffffdb514c4c51555555504c4c73ffffffffffffffffffffdb594f4c4c4c525555554f51d3ffffffffffffffffffff7b55554f4c4c4c525555554f4c4c4c525555554f4c4cdbffffffffffffffffffffc7544f4c4c4c535555544e4c4c4c5354514d4d4d5054549dffffffffffffffffffffae62656969696562626265696969656262626569696964504d4d51545454504d4d61f1ffffffffffffffffffef60504d4d4d515454545062f8fffffffffffffffffffff9eaeaeaeaeaeaeaeaeaeaeaeaeaeaeaeaeaeaeaeaeaf2ffffffffffffffffffff88544f4d4d4d525454544f6cffffffffffffffffffffdc5854544f4d4d4d52545479ffffffffffffffffffffda51525454544f4d4d4d5259d5ffffffffffffffffffff754d4d535454544e4d4d4d535454544e4d4d4d535454ddffffffffffffffffffffc54d535454544e4d4d4d535454544e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff754c4c535555554e4c4c4c535555554e4c4c4c535555ddffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff754c4c535555554e4c4c4c535555554e4c4c4c535555ddffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8955504c4c4c515555554f6bffffffffffffffffffffdc5955554f4c4c4c51555579ffffffffffffffffffffda51525555554f4c4c4c5259d5ffffffffffffffffffff754c4c525555544f4c4c4c525555544f4c4c4c525555ddffffffffffffffffffffc54d525555544e4c4c4d535555544e4d50545454504d4d9affffffffffffffffffffad54504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545468f1ffffffffffffffffffee5951545454504d4d4d5168f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff834d525454544f4d4d4d5272ffffffffffffffffffffdb514d4d525454544f4d4d73ffffffffffffffffffffdc584f4d4d4d525454544f52d4ffffffffffffffffffff7b54544e4d4d4d535454544e4d4d4d535454544e4d4ddbffffffffffffffffffffc7544e4d4d4d535454544e4d4d4d534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555568f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff834c51555555504c4c4c5172ffffffffffffffffffffdb514c4c515555554f4c4c73ffffffffffffffffffffdb594f4c4c4c525555544f51d3ffffffffffffffffffff7b55544f4c4c4c525555544f4c4c4c525555544f4c4cdbffffffffffffffffffffc7544f4c4c4d535555544e4c4c4d5354514d4d4d5054549dffffffffffffffffffffa94d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d61f1ffffffffffffffffffef60504d4d4d515454545062f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff88544f4d4d4d525454544f6cffffffffffffffffffffdc5854544f4d4d4d52545479ffffffffffffffffffffda51525454544f4d4d4d5259d5ffffffffffffffffffff754d4d535454544e4d4d4d535454544e4d4d4d535454ddffffffffffffffffffffc54d535454544e4d4d4d535454544e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff754c4c535555554e4c4c4c535555554e4c4c4c535555ddffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8fffffffffffffffffffff3f1f1f1f0f0f0f1f1f1f1f1f0f0f0f1f1f1f1f1f0f0fdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff754c4c535555554e4c4c4c535555554e4c4c4c535555ddffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffffa76d6d686666666a6d6d6d686666666a6d6d6d686666c9ffffffffffffffffffff8955504c4c4c515555554f6bffffffffffffffffffffdc5955554f4c4c4c51555579ffffffffffffffffffffda51525555554f4c4c4c5259d5ffffffffffffffffffff754c4c525555544f4c4c4c525555544f4c4c4c525555ddffffffffffffffffffffc54d525555544e4c4c4d535555544e4c50555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555568f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff834c515555554f4c4c4c5272ffffffffffffffffffffdb514c4c525555544f4c4c73ffffffffffffffffffffdc584f4c4c4c525555544f51d3ffffffffffffffffffff7b55544f4c4c4d525555544f4c4c4d525555544f4c4cdbffffffffffffffffffffc7544f4c4c4d535555544e4c4c4d534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555568f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff834c51555555504c4c4c5172ffffffffffffffffffffdb514c4c515555554f4c4c73ffffffffffffffffffffdb594f4c4c4c525555544f51d3ffffffffffffffffffff7b55544f4c4c4c525555544f4c4c4c525555544f4c4cdbffffffffffffffffffffc7544f4c4c4d535555544e4c4c4d5355514c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c61f1ffffffffffffffffffef61504c4c4c515555555062f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbeffffffffffffffffffff89554f4c4c4c515555554f6bffffffffffffffffffffdc5955544f4c4c4c52555579ffffffffffffffffffffda51525555544f4c4c4d5259d5ffffffffffffffffffff754c4d525555544f4c4c4d525555544f4c4c4d525555ddffffffffffffffffffffc54d525555544e4c4c4d535555544e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff754c4c535555554e4c4c4c535555554e4c4c4c535555ddffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff754c4c535555554e4c4c4c535555554e4c4c4c535555ddffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbeffffffffffffffffffff8955504c4c4c515555554f6bffffffffffffffffffffdc5955554f4c4c4c51555579ffffffffffffffffffffda51525555554f4c4c4c5259d5ffffffffffffffffffff754c4c525555544f4c4c4c525555544f4c4c4c525555ddffffffffffffffffffffc54d525555544e4c4c4d535555544e4c50555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555568f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff834c51555555504c4c4c5172ffffffffffffffffffffdb514c4c515555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555544f51d3ffffffffffffffffffff7b55544f4c4c4c525555544f4c4c4c525555544f4c4cdbffffffffffffffffffffc7544f4c4c4d535555544e4c4c4d534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555568f2ffffffffffffffffffee5950555555504c4c4c5069f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff834c51555555504c4c4c5172ffffffffffffffffffffdb514c4c51555554504c4c73ffffffffffffffffffffdb584f4c4c4c525555544f51d3ffffffffffffffffffff7b55544f4c4c4d525555544f4c4c4d525555544f4c4cdbffffffffffffffffffffc7544f4c4c4d535555544e4c4c4d5355514c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbeffffffffffffffffffff8955504c4c4c515555554f6bffffffffffffffffffffdc5955554f4c4c4c5155557affffffffffffffffffffda51525555554f4c4c4c5259d5ffffffffffffffffffff754c4c525555544f4c4c4c525555544f4c4c4c525555ddffffffffffffffffffffc54d525555544e4c4c4d535555544e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff754c4c535555554e4c4c4c535555554e4c4c4c535555ddffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffff754c4c535555554e4c4c4c535555554e4c4c4c535555ddffffffffffffffffffffc44c535555554e4c4c4c535555554e55514c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c505555555062f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbeffffffffffffffffffff8855504c4c4c51555555506bffffffffffffffffffffdc595554504c4c4c51555579ffffffffffffffffffffda51525555544f4c4c4d5259d5ffffffffffffffffffff754c4d525555544f4c4c4d525555544f4c4c4d525555ddffffffffffffffffffffc54d525555544e4c4c4d535555544e4c50555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555568f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff834c51555555504c4c4c5172ffffffffffffffffffffdb514c4c515555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555544f51d3ffffffffffffffffffff7b55544f4c4c4c525555544f4c4c4c525555544f4c4cdbffffffffffffffffffffc7544f4c4c4d535555544e4c4c4d534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffff7c55554e4c4c4c535555554e4c4c4c535555554e4c4cdbffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534d4f545454514d4d99ffffffffffffffffffffac54514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545468f2ffffffffffffffffffee5a50545454514d4d4d5068f8ffffffffffffffffffff954d4d50545454504d4d4d51545454504d4d4d515454c0ffffffffffffffffffff834d51545454504d4d4d5172ffffffffffffffffffffdb514d4d51545454504d4d73ffffffffffffffffffffdb58504d4d4d515454545052d3ffffffffffffffffffff7b54544f4d4d4d525454544f4d4d4d525454544f4d4ddbffffffffffffffffffffc7544f4d4d4d525454544f4d4d4d5255514c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbeffffffffffffffffffff8955504c4c4c515555554f6bffffffffffffffffffffdc5955554f4c4c4c5155557affffffffffffffffffffda51525555554f4c4c4c5259d5ffffffffffffffffffff754c4c525555544f4c4c4c525555544f4c4c4c525555ddffffffffffffffffffffc54d525555544e4c4c4d535555544e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffffc1aaaaacaeaeaeabaaaaaaacaeaeaeabaaaaaaacaeaeecffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc44c535555554e4c4c4c535555554e54524d4d4d4f54549effffffffffffffffffffaa4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d61f1ffffffffffffffffffee60514d4d4d505454545162f8ffffffffffffffffffff995454504d4d4d51545454504d4d4d51545454504d4dbeffffffffffffffffffff8854504d4d4d51545454506cffffffffffffffffffffdc585454504d4d4d51545479ffffffffffffffffffffda5151545454504d4d4d5159d5ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc54d525454544f4d4d4d525454544f4c50555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555568f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff834c51555555504c4c4c5172ffffffffffffffffffffdb514c4c515555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555544f51d3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7544f4c4c4d535555544e4c4c4d534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534c4f555555514c4c99ffffffffffffffffffffad55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555569f2ffffffffffffffffffee5951555555504c4c4c5169f8ffffffffffffffffffff954c4c51555555504c4c4c51555555504c4c4c515555c0ffffffffffffffffffff824c525555554f4c4c4c5273ffffffffffffffffffffdb504c4c525555554f4c4c73ffffffffffffffffffffdc594f4c4c4c525555554f51d3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7554e4c4c4c535555554e4c4c4c534d4f545454514d4d99ffffffffffffffffffffac54514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545468f2ffffffffffffffffffee5a50545454514d4d4d5068f8ffffffffffffffffffff954d4d50545454504d4d4d51545454504d4d4d515454c0ffffffffffffffffffff834d51545454504d4d4d5172ffffffffffffffffffffdb514d4d51545454504d4d73ffffffffffffffffffffdb58504d4d4d515454545052d3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7544f4d4d4d525454544f4d4d4d5255514c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c505555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbeffffffffffffffffffff89554f4c4c4c515555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda51525555554f4c4c4c5259d5ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc54c525555544e4c4c4c535555544e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc44c535555554e4c4c4c535555554e55524c4c4c5055559effffffffffffffffffffa94c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c61f1ffffffffffffffffffef61504c4c4c515555555061f8ffffffffffffffffffff9a5555504c4c4c51555555504c4c4c51555555504c4cbdffffffffffffffffffff89554f4c4c4c525555554f6bffffffffffffffffffffdc5955554f4c4c4c5255557affffffffffffffffffffda50525555554f4c4c4c525ad5ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc44c535555554e4c4c4c535555554e54524d4d4d5054549effffffffffffffffffffaa4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d61f1ffffffffffffffffffee60514d4d4d505454545162f8ffffffffffffffffffff995454504d4d4d51545454504d4d4d51545454504d4dbeffffffffffffffffffff8854504d4d4d51545454506cffffffffffffffffffffdc585454504d4d4d51545479ffffffffffffffffffffda5151545454504d4d4d5159d5ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc54d525454544f4d4d4d525454544f4c4f555555514c4c6fa4a7a7a7a4a2a2a2a4a78155514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c505555609ba2a2a2a4a7a7a7a4a2995350555555504c4c4c5060a4a7a4a2a2a2a4a7a7a7a46f4c4c51555555504c4c4c51555555504c4c4c51555588a4a2a2a2a5a7a7a7a3a2694c515555554f4c4c4c5262a7a7a3a2a2a2a5a7a7a7934f4c4c525555554f4c4c61a5a7a7a7a3a2a2a2a5a797574f4c4c4c525555554f4f8aa2a5a7a7a6a3a2a2a2a5a7a7a6a3a2a2a2a5a7a7a6a3a2a2a2a5a7a7a6a3a2a2a2a5a7a7a6a3a2a2a2a5a78d544f4c4c4c535555544e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534d4f545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d515454544f4d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4d4d4d5255514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c515555554f4c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555544f4c4c4c525555544f4c4c4c525555544e4c4c4c535555544e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e54514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555544f4c4c4c525555544f4c4c4c535555544e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534d50545454514d4d3e2d2f2f2f2e2b2b2b2d2f2f2f2e2b2b2b2d2f2f2f2e2b2b2b2d2f2f2f2e2b2b2b2d2f2f2f2d2b2b2b2d2f2f2f2d2b2b2b2d2f2f2f2d2b2f4b50545454514d4d4d5050322f2d2b2b2b2e2f2f2f2d404d4d51545454504d4d4d3b2f2f2f2d2b2b2b2e2f2f46504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454492c2b2b2e2f2f2f2d2b2b2b2e2f2f2f2d2b2b2b2e2f2f2f2d2b2b2b2e2f2f2f2d2c474d51545454504d4d4d51382f2f2c2b2b2b2e2f2f2f2c2b2b2b2e2f2f2f2c2b2b2b2e2f2f2f2c2b2b2b2e2f3b544f4d4d4d525454544f4d4d4d5255514c4c4c505555391515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151b50504c4c4c50555555504617151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c515555554f4c4c4c515555554f4c4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c525555544e4c4c4c535555544e55524c4c4c505555391515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151b50504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c535555554e4c4c4c535555554e55524c4c4c505555391515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151b50504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c535555554e4c4c4c535555554e54514d4d4d505454391515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151b4f514d4d4d50545454514717151515151515151515153a5454504d4d4d515454542c151515151515151515153951545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d441615151515151515151515151515151515151515151515151515151515151515174454504d4d4d5154545450221515151515151515151515151515151515151515151515151515151515151515284d525454544f4d4d4d525454544f4c50555555514c4c341515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151a4851555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153d504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151515151515151515151515151515151515151515151515163f4c525555554f4c4c4c522315151515151515151515151515151515151515151515151515151515151515152a554e4c4c4c535555554e4c4c4c534c4f555555514c4c341515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151a4851555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151515151515151515151515151515151515151515151515163f4c525555554f4c4c4c522315151515151515151515151515151515151515151515151515151515151515152a554e4c4c4c535555554e4c4c4c534c4f555555514c4c341515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151a4851555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151515151515151515151515151515151515151515151515163f4c525555554f4c4c4c522315151515151515151515151515151515151515151515151515151515151515152a554e4c4c4c535555554e4c4c4c534d4f545454514d4d351515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151b4a50545454514d4d4d504c1715151515151515151515374d4d51545454504d4d4d2a151515151515151515153c504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d5154545345161515151515151515151515151515151515151515151515151515151515151517404d51545454504d4d4d5123151515151515151515151515151515151515151515151515151515151515151529534f4d4d4d525454534f4d4d4d5255514c4c4c505555391515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151b50504c4c4c51555555504617151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c525555554e4c4c4c535555554e55524c4c4c505555391515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151515151b50504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c535555554e4c4c4c535555554e55524c4c4c5055553e1e1d1d1d1e1f1f1f1e1d1d1d1e1f1f1f1e1d1d1d1e1e15151515151515151515151d1d1d1e1f1f1f1e1d1d1d1e1f1f1f1e1d1d1d1e1f2451504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515171e1d1d1d1f1f1f1f1e1d1d1d1f1f1f1f1e1d1d1d1f2047554f4c4c4c525555554f22151515151515151515151d1f1f1f1e1d1d1d1f1f1f1f1e1d1d1d1f1f1f1f1e1d2c4c535555554e4c4c4c535555554e54514d4d4d505454544f4b4b4b4e5151514f4b4b4b4e5151514f4b4b4b4e4c1915151515151515151518484b4b4e5151514e4b4b4b4e5151514e4b4b4b4e515153514d4d4d50545454514717151515151515151515153a5454504d4d4d515454542c151515151515151515153951545454504d4d4d51545454504d4d4d51545454504d4d4d51545453504d4d4d4416151515151515151515224e4b4b4b4f5151514e4b4b4b4f5151514e4b4b4b4f515254504d4d4d51545454502215151515151515151517465151514d4b4b4b4f5151514d4b4b4b4f5151514d4b4b4d525454534f4d4d4d525454534f4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153d504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c522315151515151515151517424c4c4c525555554e4c4c4c525555554e4c4c4c525555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c522315151515151515151517424c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c522315151515151515151517424c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534e4f535353514e4e4e4f535353514e4e4e50535353514e4e4e50535353514919151515151515151515184e5353514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504c1715151515151515151515374e4e50535353504e4e4e2a151515151515151515153c504e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e5053535345161515151515151515152151535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e512315151515151515151517444e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e525353534f4e4e4e5255514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504617151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f2215151515151515151517485555554e4c4c4c525555554e4c4c4c525555554e4c4c4c525555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f2215151515151515151517485555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f2215151515151515151517485555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e53524e4e4e4f535353514e4e4e4f535353514e4e4e50535353514e4e4e504e1a151515151515151515184a4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e5053535351471715151515151515151515395353504e4e4e515353532c151515151515151515153951535353514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e441615151515151515151522504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e5153535350221515151515151515151746535353504e4e4e51535353504e4e4e51535353504e4e4e515353534f4e4e4e525353534f4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153d504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c522315151515151515151517424c4c4c525555554e4c4c4c525555554e4c4c4c525555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c522315151515151515151517424c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c522315151515151515151517424c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534e4f535353514e4e4e4f535353514e4e4e50535353514e4e4e50535353514919151515151515151515184e5353514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504c1715151515151515151515374e4e50535353504e4e4e2a151515151515151515153c504e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e5053535345161515151515151515152151535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e512315151515151515151517444e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e525353534f4e4e4e5255514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504617151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f2215151515151515151517485555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f2215151515151515151517485555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f2215151515151515151517485555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e53524e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504d1a151515151515151515184a4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e5053535351471715151515151515151515395353504e4e4e515353532c151515151515151515153951535353514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e441615151515151515151522504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e5153535350221515151515151515151746535353504e4e4e51535353504e4e4e51535353504e4e4e515353534f4e4e4e515353534f4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153d504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c522315151515151515151517424c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c522315151515151515151517424c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c522315151515151515151517424c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534e4f535353514e4e4e50535353514e4e4e50535353514e4e4e50535353514919151515151515151515184e5353514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504c1715151515151515151515374e4e51535353504e4e4e2a151515151515151515153c504e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e5053535345161515151515151515152151535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e512315151515151515151517444e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e515353534f4e4e4e5155514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504617151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c45161515151515151515152045434343474a4a4a45434343474a4a4a45434343474a54554f4c4c4c525555554f22151515151515151515163e4a4a4a45434343484a4a4a45434343484a4a4a4543464c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c535555554e4c4c4c535555554e53514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504d1a151515151515151515184a4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e5053535351481715151515151515151515395353504e4e4e515353532c151515151515151515153951535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e441615151515151515151515151515151515151515151515151515151515151515174353504e4e4e5153535350221515151515151515151515151515151515151515151515151515151515151515284e515353534f4e4e4e525353534f4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153d504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151515151515151515151515151515151515151515151515163f4c525555554f4c4c4c522315151515151515151515151515151515151515151515151515151515151515152a554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151515151515151515151515151515151515151515151515163f4c525555554f4c4c4c522315151515151515151515151515151515151515151515151515151515151515152a554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151515151515151515151515151515151515151515151515163f4c525555554f4c4c4c522315151515151515151515151515151515151515151515151515151515151515152a554e4c4c4c535555554e4c4c4c534e50535353514e4e4e50535353514e4e4e50535353514e4e4e50535353514919151515151515151515184e5353514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504b1715151515151515151515374e4e51535353504e4e4e2a151515151515151515153c504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e5153535345161515151515151515151515151515151515151515151515151515151515151517404e51535353504e4e4e5123151515151515151515151515151515151515151515151515151515151515151529534f4e4e4e525353534f4e4e4e5255514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504617151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c535555554e4c4c4c535555554e53514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504d1a151515151515151515184a4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e5053535351481715151515151515151515395353504e4e4e515353532c151515151515151515153951535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e441615151515151515151517212121212020202021212121202020202121212120214653504e4e4e51535353502c2121202020202121212120202020212121212020201715151515151515151515284e515353534f4e4e4e525353534f4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521505353534d4b4b4b505353534d4b4b4b515353534d4b4c4c525555554f4c4c4c525453534d4b4b4b515353534d4b4b4b515353534d4b4b20151515151515151515152a554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c20151515151515151515152a554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c20151515151515151515152a554e4c4c4c535555554e4c4c4c534e50535353514e4e4e50535353514e4e4e50535353514e4e4e50535353514919151515151515151515184e5353504e4e4e50535353504e4e4e50535353514e4e4e50535353504e4e4e504b1715151515151515151515374e4e51535353504e4e4e2a151515151515151515153c504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e5153535245161515151515151515152151535352504e4e4e51535352504e4e4e51535353504e4e4e51535353504e4e4e515353534f4e4e4e515353534f4e4e4e51535353504e4e20151515151515151515152952504e4e4e525353524f4e4e4e5255514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504617151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c5355552215151515151515151515274c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c5355552215151515151515151515274c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c5355552215151515151515151515274c535555554e4c4c4c535555554e53514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504d1a151515151515151515184a4e4e50535353504e4e4e50535353514e4e4e50535353504e4e4e5053535350481715151515151515151515395353504e4e4e515353532c151515151515151515153951535353504e4e4e51535353504e4e4e51535353504e4e4e51535352504e4e4e441615151515151515151522504e4e4e51535352504e4e4e51535352504e4e4e51535353504e4e4e51535353504e4e4e515353534f4e4e4e51535353504e4e4e5153532115151515151515151515284e515353524f4e4e4e525353524f4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c20151515151515151515152a554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c20151515151515151515152a554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c20151515151515151515152a554e4c4c4c535555554e4c4c4c534f4f525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514919151515151515151515184e5252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f504b1715151515151515151515384f4f50525252514f4f4f2a151515151515151515153b504f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f5052525245161515151515151515152251525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f20151515151515151515152852504f4f4f51525252504f4f4f5155514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504617151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c5355552215151515151515151515274c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c5355552215151515151515151515274c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c5355552215151515151515151515274c535555554e4c4c4c535555554e52524f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f504d1a151515151515151515184b4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f5052525251481715151515151515151515395252504f4f4f505252522c151515151515151515153a50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f441615151515151515151522504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f5152522115151515151515151515284f51525252504f4f4f51525252504c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c20151515151515151515152a554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c20151515151515151515152a554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a151515151515151515153e504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555441615151515151515151521525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c20151515151515151515152a554e4c4c4c535555554e4c4c4c534f4f525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514919151515151515151515184e5252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f504b1715151515151515151515384f4f50525252514f4f4f2a151515151515151515153b504f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f5052525245161515151515151515152251525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f20151515151515151515152852504f4f4f51525252504f4f4f5155514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c5355552215151515151515151515274c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c1515151515151515151538515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c4516151515151515151515234f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c5355552215151515151515151515274c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c151515151515151515151d2425252524222222242525252422222224252525242a4c4c525555554f4c4c4c451615151515151515151518242222232425252524222223242525252422222324264b554f4c4c4c525555554f2c2223242525252322222324252525232222232425251815151515151515151515274c535555554e4c4c4c535555554e52524f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f504d1a151515151515151515184b4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f5052525251481715151515151515151515395252514f4f4f505252522c15151515151515151515151515151515151515151515151515151515151515151f4f4f50525252514f4f4f441615151515151515151515151515151515151515151515151515151515151515174352504f4f4f5152525250221515151515151515151515151515151515151515151515151515151515151515284f51525252504f4f4f51525252504c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a15151515151515151515151515151515151515151515151515151515151515152055554f4c4c4c52555555441615151515151515151515151515151515151515151515151515151515151515163f4c525555554f4c4c4c522315151515151515151515151515151515151515151515151515151515151515152a554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a15151515151515151515151515151515151515151515151515151515151515152055554f4c4c4c52555555441615151515151515151515151515151515151515151515151515151515151515163f4c525555554f4c4c4c522315151515151515151515151515151515151515151515151515151515151515152a554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471915151515151515151518505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514d1715151515151515151515364c4c51555555504c4c4c2a15151515151515151515151515151515151515151515151515151515151515152055554f4c4c4c52555555441615151515151515151515151515151515151515151515151515151515151515163f4c525555554f4c4c4c522315151515151515151515151515151515151515151515151515151515151515152a554e4c4c4c535555554e4c4c4c534f4f525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514a19151515151515151515184d5252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f504b1715151515151515151515384f4f50525252514f4f4f2a15151515151515151515151515151515151515151515151515151515151515151f5252514f4f4f5052525245161515151515151515151515151515151515151515151515151515151515151517414f51525252504f4f4f512315151515151515151515151515151515151515151515151515151515151515152852504f4f4f51525252504f4f4f5155514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c15151515151515151515151515151515151515151515151515151515151515151f4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c15151515151515151515151515151515151515151515151515151515151515151f4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1a15151515151515151518484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504517151515151515151515153b5555504c4c4c515555552c15151515151515151515151515151515151515151515151515151515151515151f4c4c525555554f4c4c4c4516151515151515151515151515151515151515151515151515151515151515151745554f4c4c4c525555554f221515151515151515151515151515151515151515151515151515151515151515274c535555554e4c4c4c535555554e52514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f504c1a151515151515151515184b4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f5052525251481715151515151515151515395252504f4f4f515252522b15151515151515151515151515151515151515151515151515151515151515151f4f4f50525252504f4f4f441615151515151515151515151515151515151515151515151515151515151515174252514f4f4f5052525251221515151515151515151515151515151515151515151515151515151515151515284f51525252504f4f4f51525252504c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471b1717171717171717171a505555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c514e1a17171717171717171717364c4c51555555504c4c4c2b17171717171717171717171717171717171717171717171717171717171717172155554f4c4c4c52555555451817171717171717171717171717171717171717171717171717171717171717183f4c525555554f4c4c4c522517171717171717171717171717171717171717171717171717171717171717172b554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4240434747474340404043535555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51544747434040404447474743464c4c51555555504c4c4c4947474743404040444747474340404044474747424040404447474742404040444855554f4c4c4c525555554f404040444747474240404045474747424040404547474742404040454747474240474c525555554f4c4c4c524a47474240404045474747424040404547474742404040454747474240404045474a554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f50525252514f4f4f50525252514f4f4f50525252504f4f4f50525252504f4f4f50525252504f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f5155524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e52514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252514f4f4f50525252514f4f4f50525252504f4f4f50525252504f4f4f50525252504f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525251514f4f4f50525251514f4f4f50525251514f4f4f50525251514f4f4f50525252514f4f4f50525252514f4f4f50525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f5155524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e;
parameter [88451:0] ROM_G = 88452'h4c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c5353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e515353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c515555554f4c4c4c515555554f4c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c525555554e4c4c4c525555554e4c4c4c525555554e4c4c4c535555554e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e525353534f4e4e4e524c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c50555959595653535355595959565353535559595956535353555959595653535355555555514c4c4c5055555556535353555959595653524c51555555504c4c4c515559595553535356595959555353535659595955535353565959595553535356595959555353535659595955534d4c525555554f4c4c4c5256595955535353565959595553535356595959555353535659595955535353565958554f4c4c4c525555554f4c525356595959555353535659595954535353575959595453535357595959545353535759595954535353575957554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161616161616161616161616161616161616161616161616160565555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51566161616161616161616161616161616161616161616161616161616161616161616161616161616161616161534c51555555504c4c4c515761616161616161616161616161616161616161616161616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161616161616161616161616161616161616161616161616161616161616161616161615d554e4c4c4c535555554e4c4c4c5353504e4e4e515353596161616161616161616161616161616161616161616161616161616161616161604f4e4e51535353504e4e50606161616161616161616054504e4e4e515353535050606161616161616161616161616161616161616161616161616161616161616161616161616161616161616158534f4e4e4e525353534f5161616161616161616161616161616161616161616161616161616161616161615d4e525353534f4e4e4e52535d616161616161616161616161616161616161616161616161616161616161616161616161616161616161615a4e525353534f4e4e4e525353534f55524c4c4c5055555a6161616161616161616161616161616161616161616161616161616161616161604e4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e606161616161616161616161616161616161616161616161616161616161616161616161616161616161616159554f4c4c4c525555554f4f61616161616161616161616161616161616161616161616161616161616161615d4d525555554f4c4c4c52555e616161616161616161616161616161616161616161616161616161616161616161616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a6161616161616161616161616161616161616161616161616161616161616161604e4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e606161616161616161616161616161616161616161616161616161616161616161616161616161616161616159554f4c4c4c525555554f4f61616161616161616161616161616161616161616161616161616161616161615d4d525555554f4c4c4c52555e616161616161616161616161616161616161616161616161616161616161616161616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a6161616161616161616161616161616161616161616161616161616161616161604e4c4c50555555514c4c4f5f6161616161616161616056504c4c4c51555555504f60616161616161616161616161616161616161616161616161616161616161616161616161616161616161615855504c4c4c515555554f5061616161616161616161616161616161616161616161616161616161616161615d4d525555554f4c4c4c52555e616161616161616161616161616161616161616161616161616161616161616161616161616161616161615a4c525555554e4c4c4c535555554e4d50545454504d4d56616161616161616161616161616161616161616161616161616161616161616160555454504d4d4d51545455606161616161616161615f4f51545454504d4d4d51556061616161616161616161616161616161616161616161616161616161616161616161616161616161616161534d515454544f4d4d4d525661616161616161616161616161616161616161616161616161616161616161615e544f4d4d4d525454534f4e5c616161616161616161616161616161616161616161616161616161616161616161616161616161616161615d534f4d4d4e535454534e4d4d4e534c4f555555514c4c55616161616161616161616161616161616161616161616161616161616161616160565555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161616161616161616161616161616161616161616161616161616161616161616161524c525555554f4c4c4c525761616161616161616161616161616161616161616161616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161616161616161616161616161616161616161616161616161616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161616161616161616161616161616161616161616161616160565555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161616161616161616161616161616161616161616161616161616161616161616161524c525555554f4c4c4c525761616161616161616161616161616161616161616161616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161616161616161616161616161616161616161616161616161616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161616161616161616161616161616161616161616161616160565555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51566161616161616161616161616161616161616161616161616161616161616161616161616161616161616161534c51555555504c4c4c515761616161616161616161616161616161616161616161616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161616161616161616161616161616161616161616161616161616161616161616161615d554e4c4c4c535555554e4c4c4c5354514d4d4d515454596161616161616161616161616161616161616161616161616161616161616161604f4d4d51545454504d4d50606161616161616161616055504d4d4d515454545050606161616161616161616161616161616161616161616161616161616161616161616161616161616161616158544f4d4d4d515454544f5161616161616161616161616161616161616161616161616161616161616161615d4e525454534f4d4d4e52545e616161616161616161616161616161616161616161616161616161616161616161616161616161616161615a4e525454534e4d4d4e535454534e55524c4c4c5055555a6161616161616161616161616161616161616161616161616161616161616161604e4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e606161616161616161616161616161616161616161616161616161616161616161616161616161616161616159554f4c4c4c525555554f4f61616161616161616161616161616161616161616161616161616161616161615d4d525555554f4c4c4c52555e616161616161616161616161616161616161616161616161616161616161616161616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a6161616161616161616158505357575753505050535860616161616161616161604e4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615b5757535050505457575753505050545757575350505b6161616161616161616159554f4c4c4c525555554f4f616161616161616161615f5757575250505054575759616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161545050555757575150505055575757515050505557575f616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c505660616161616161616161604e4c4c50555555514c4c4f5f6161616161616161616056504c4c4c51555555504f60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c59616161616161616161615855504c4c4c515555554f50616161616161616161615e5555554f4c4c4c51555557616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c525555554f4c4c4c525555554e4c4c4c5255555f616161616161616161615a4c525555554e4c4c4c535555554e4d50545454504d4d56616161616161616161615b54504d4d4d51545454504f6061616161616161616160555454504d4d4d51545455606161616161616161615f4f51545454504d4d4d51556161616161616161616161554d4d51545454504d4d4d51545454504d4d4d5154545c61616161616161616161534d51545454504d4d4d5156616161616161616161615d4e4d4d515454544f4d4d52616161616161616161615e544f4d4d4d525454534f4e5c616161616161616161615754534f4d4d4d525454534f4d4d4d525454534f4d4d5d616161616161616161615d534f4d4d4e535454534e4d4d4e534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514e5f61616161616161616160565555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514e5f61616161616161616160565555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514e5f61616161616161616160565555514c4c4c50555556606161616161616161615f4e50555555504c4c4c50566161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555c61616161616161616161534c51555555504c4c4c5157616161616161616161615d4d4c4c51555555504c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554f4c4c4c525555554f4c4c4c525555554f4c4c5d616161616161616161615d544f4c4c4c535555544e4c4c4c5354514d4d4d5154545961616161616161616161574d51545454504d4d4d515560616161616161616161604f4d4d51545454504d4d50606161616161616161616055504d4d4d5154545450506061616161616161616161595454504d4d4d51545454504d4d4d51545454504d4d5a616161616161616161615854504d4d4d515454544f51616161616161616161615e5454544f4d4d4d51545456616161616161616161615d4e525454544f4d4d4d52545e61616161616161616161524d4d525454534f4d4d4d525454534f4d4d4d5254545e616161616161616161615a4e525454534e4d4d4e535454534e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c505660616161616161616161604e4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c535555554e4c4c4c535555554e4c4c4c5355555f616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c505660616161616161616161604e4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c535555554e4c4c4c535555554e4c4c4c5355555f616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c505660616161616161616161604e4c4c50555555514c4c4f5f6161616161616161616056504c4c4c50555555504f60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c59616161616161616161615855504c4c4c515555555050616161616161616161615e555555504c4c4c51555557616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c525555554f4c4c4c525555554f4c4c4c5255555f616161616161616161615a4c525555544e4c4c4c535555544e4d50545454504d4d56616161616161616161615b54514e4e4e5254545451506061616161616161616160555454504d4d4d51545455606161616161616161615f4f51545454504d4d4d51556161616161616161616161554d4d51545454504d4d4d51545454504d4d4d5154545c61616161616161616161534d51545454504d4d4d5156616161616161616161615d4e4d4d515454544f4d4d52616161616161616161615e544f4d4d4d525454534f4e5c616161616161616161615754534f4d4d4d525454534f4d4d4d525454534f4d4d5d616161616161616161615d534f4d4d4e535454534e4d4d4e534c4f555555514c4c5561616161616161616161605f5e5d5d5d5e5f5f5f5e5e6161616161616161616160565555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161616161616161616161616161616161616161616161616160565555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161616161616161616161616161616161616161616161616160565555514c4c4c50555556606161616161616161615f4e50555555504c4c4c50566161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555c61616161616161616161534c51555555504c4c4c5157616161616161616161615d4d4c4c51555555504c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554f4c4c4c525555554f4c4c4c525555554f4c4c5d616161616161616161615d544f4c4c4c535555544e4c4c4c5354514d4d4d505454596161616161616161616161616161616161616161616161616161616161616161604e4d4d51545454504d4d4f606161616161616161616055504d4d4d51545454504f6061616161616161616161595454504d4d4d51545454504d4d4d51545454504d4d5a6161616161616161616158544f4d4d4d525454544f50616161616161616161615e5454544f4d4d4d52545457616161616161616161615d4d525454544f4d4d4d52545e61616161616161616161524d4d535454544e4d4d4d535454544e4d4d4d5354545e616161616161616161615a4d535454544e4d4d4d535454544e55524c4c4c5055555a6161616161616161616161616161616161616161616161616161616161616161604e4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c535555554e4c4c4c535555554e4c4c4c5355555f616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a6161616161616161616161616161616161616161616161616161616161616161604e4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c535555554e4c4c4c535555554e4c4c4c5355555f616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a6161616161616161616161616161616161616161616161616161616161616161604e4c4c50555555514c4c4f5f6161616161616161616056504c4c4c50555555504f60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c59616161616161616161615855504c4c4c515555555050616161616161616161615e555555504c4c4c51555557616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c525555554f4c4c4c525555554f4c4c4c5255555f616161616161616161615a4c525555544e4c4c4c535555544e4d50545454514d4d56616161616161616161616161616161616161616161616161616161616161616160555454504d4d4d51545455606161616161616161615f4e51545454504d4d4d51566161616161616161616161554d4d51545454504d4d4d51545454504d4d4d5154545c61616161616161616161534d525454544f4d4d4d5256616161616161616161615d4d4d4d525454544f4d4d51616161616161616161615e544f4d4d4d525454544f4d5c616161616161616161615754544e4d4d4d535454544e4d4d4d535454544e4d4d5d616161616161616161615d544e4d4d4d535454544e4d4d4d534c4f555555514c4c55616161616161616161616161616161616161616161616161616161616161616160565555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161616161616161616161616161616161616161616161616160565555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161616161616161616161616161616161616161616161616160565555514c4c4c50555556606161616161616161615f4e50555555504c4c4c50566161616161616161616161554d4d51555555504d4d4d51555555504d4d4d5155555d61616161616161616161534c51555555504c4c4c5157616161616161616161615d4d4c4c51555555504c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554f4c4c4c525555554f4c4c4c525555554f4c4c5d616161616161616161615d544f4c4c4c535555544e4c4c4c5354514d4d4d5054545961616161616161616161584f52565656524f4f4f52565656524f4f4f52565656524d4d4d51545454504d4d4f606161616161616161616055504d4d4d51545454504f6061616161616161616161615f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f5f606161616161616161616158544f4d4d4d525454544f50616161616161616161615e5454544f4d4d4d52545457616161616161616161615d4d525454544f4d4d4d52545e61616161616161616161514d4d535454544e4d4d4d535454544e4d4d4d5354545e616161616161616161615a4d535454544e4d4d4d535454544e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e606161616161616161616161616161616161616161616161616161616161616161616161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c535555554e4c4c4c535555554e4c4c4c5355555f616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e606161616161616161616161616161616161616161616161616161616161616161616161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c535555554e4c4c4c535555554e4c4c4c5355555f616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4f5f6161616161616161616056504c4c4c51555555504f60616161616161616161616161616161616161616161616161616161616161616161616161616161616161615855504c4c4c515555554f50616161616161616161615e5555554f4c4c4c51555557616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c525555544f4c4c4c525555544f4c4c4c5255555f616161616161616161615a4d525555544e4c4c4d535555544e4d50545454504d4d56616161616161616161615b54504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545455606161616161616161615f4e51545454504d4d4d51566161616161616161616161616161616161616161616161616161616161616161616161616161616161616161534d525454544f4d4d4d5256616161616161616161615d4d4d4d525454544f4d4d51616161616161616161615e544f4d4d4d525454544f4d5c616161616161616161615754544e4d4d4d535454544e4d4d4d535454544e4d4d5d616161616161616161615d544e4d4d4d535454544e4d4d4d534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161616161616161616161616161616161616161616161616161616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161616161616161616161616161616161616161616161616161616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51566161616161616161616161616161616161616161616161616161616161616161616161616161616161616161534c51555555504c4c4c5157616161616161616161615d4d4c4c515555554f4c4c51616161616161616161615e554f4c4c4c525555544f4d5c616161616161616161615855544f4c4c4c525555544f4c4c4c525555544f4c4c5d616161616161616161615d544f4c4c4d535555544e4c4c4d5354514d4d4d5054545961616161616161616161574d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4f606161616161616161616055504d4d4d51545454504f606161616161616161616161616161616161616161616161616161616161616161616161616161616161616158544f4d4d4d525454544f50616161616161616161615e5454544f4d4d4d52545457616161616161616161615d4d525454544f4d4d4d52545e61616161616161616161514d4d535454544e4d4d4d535454544e4d4d4d5354545e616161616161616161615a4d535454544e4d4d4d535454544e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e606161616161616161616161616161616161616161616161616161616161616161616161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c535555554e4c4c4c535555554e4c4c4c5355555f616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161616060605f5f5f5f606060605f5f5f5f606060605f5f5f616161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c535555554e4c4c4c535555554e4c4c4c5355555f616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4f5f6161616161616161616056504c4c4c51555555504f60616161616161616161615a5656524f4f4f53565656524f4f4f53565656524f4f5b616161616161616161615855504c4c4c515555554f50616161616161616161615e5555554f4c4c4c51555557616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c525555544f4c4c4c525555544f4c4c4c5255555f616161616161616161615a4d525555544e4c4c4d535555544e4c50555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555556606161616161616161615f4e51555555504c4c4c51566161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555c61616161616161616161534c515555554f4c4c4c5257616161616161616161615d4d4c4c525555544f4c4c51616161616161616161615e554f4c4c4c525555544f4d5c616161616161616161615755544f4c4c4d525555544f4c4c4d525555544f4c4c5d616161616161616161615d544f4c4c4d535555544e4c4c4d534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51566161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555c61616161616161616161534c51555555504c4c4c5157616161616161616161615d4d4c4c515555554f4c4c51616161616161616161615e554f4c4c4c525555544f4d5c616161616161616161615855544f4c4c4c525555544f4c4c4c525555544f4c4c5d616161616161616161615d544f4c4c4d535555544e4c4c4d5355514c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4f5f6161616161616161616055504c4c4c51555555504f60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616158554f4c4c4c515555554f50616161616161616161615e5555544f4c4c4c52555557616161616161616161615d4d525555544f4c4c4d52555e61616161616161616161514c4d525555544f4c4c4d525555544f4c4c4d5255555f616161616161616161615a4d525555544e4c4c4d535555544e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c535555554e4c4c4c535555554e4c4c4c5355555f616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c535555554e4c4c4c535555554e4c4c4c5355555f616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4f5f6161616161616161616056504c4c4c51555555504f60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c59616161616161616161615855504c4c4c515555554f50616161616161616161615e5555554f4c4c4c51555557616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c525555544f4c4c4c525555544f4c4c4c5255555f616161616161616161615a4d525555544e4c4c4d535555544e4c50555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51566161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555c61616161616161616161534c51555555504c4c4c5157616161616161616161615d4d4c4c515555554f4c4c51616161616161616161615e554f4c4c4c525555544f4d5c616161616161616161615855544f4c4c4c525555544f4c4c4c525555544f4c4c5d616161616161616161615d544f4c4c4d535555544e4c4c4d534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e50555555504c4c4c50566161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555c61616161616161616161534c51555555504c4c4c5157616161616161616161615d4d4c4c51555554504c4c51616161616161616161615e554f4c4c4c525555544f4d5c616161616161616161615755544f4c4c4d525555544f4c4c4d525555544f4c4c5d616161616161616161615d544f4c4c4d535555544e4c4c4d5355514c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4f5f6161616161616161616056504c4c4c51555555504f60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c59616161616161616161615855504c4c4c515555554f50616161616161616161615e5555554f4c4c4c51555557616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c525555544f4c4c4c525555544f4c4c4c5255555f616161616161616161615a4d525555544e4c4c4d535555544e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c535555554e4c4c4c535555554e4c4c4c5355555f616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c535555554e4c4c4c535555554e4c4c4c5355555f616161616161616161615a4c535555554e4c4c4c535555554e55514c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4f5f6161616161616161616055504c4c4c50555555504f6061616161616161616161595555504c4c4c51555555504c4c4c51555555504c4c59616161616161616161615855504c4c4c515555555050616161616161616161615e555554504c4c4c51555557616161616161616161615d4d525555544f4c4c4d52555e61616161616161616161514c4d525555544f4c4c4d525555544f4c4c4d5255555f616161616161616161615a4d525555544e4c4c4d535555544e4c50555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51566161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555c61616161616161616161534c51555555504c4c4c5157616161616161616161615d4d4c4c515555554f4c4c51616161616161616161615e554f4c4c4c525555544f4d5c616161616161616161615855544f4c4c4c525555544f4c4c4c525555544f4c4c5d616161616161616161615d544f4c4c4d535555544e4c4c4d534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161615855554e4c4c4c535555554e4c4c4c535555554e4c4c5d616161616161616161615d554e4c4c4c535555554e4c4c4c534d4f545454514d4d55616161616161616161615b54514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545456606161616161616161615f4e50545454514d4d4d50566161616161616161616161554d4d50545454504d4d4d51545454504d4d4d5154545c61616161616161616161534d51545454504d4d4d5156616161616161616161615d4d4d4d51545454504d4d51616161616161616161615e54504d4d4d51545454504d5c616161616161616161615754544f4d4d4d525454544f4d4d4d525454544f4d4d5d616161616161616161615d544f4d4d4d525454544f4d4d4d5255514c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4f5f6161616161616161616056504c4c4c51555555504f60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c59616161616161616161615855504c4c4c515555554f50616161616161616161615e5555554f4c4c4c51555557616161616161616161615d4d525555554f4c4c4c52555e61616161616161616161514c4c525555544f4c4c4c525555544f4c4c4c5255555f616161616161616161615a4d525555544e4c4c4d535555544e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e616161616161616161615a57575a5b5b5b585757575a5b5b5b585757575a5b5b60616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e616161616161616161616161616161616161616161616161616161616161616161616161616161616161615a4c535555554e4c4c4c535555554e54524d4d4d4f54545a61616161616161616161584d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4f5f6161616161616161615f55514d4d4d50545454514f6061616161616161616161595454504d4d4d51545454504d4d4d51545454504d4d59616161616161616161615854504d4d4d515454545050616161616161616161615e545454504d4d4d51545457616161616161616161615d4d51545454504d4d4d51555e616161616161616161616161616161616161616161616161616161616161616161616161616161616161615a4d525454544f4d4d4d525454544f4c50555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51566161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555c61616161616161616161534c51555555504c4c4c5157616161616161616161615d4d4c4c515555554f4c4c51616161616161616161615e554f4c4c4c525555544f4d5c616161616161616161616161616161616161616161616161616161616161616161616161616161616161615d544f4c4c4d535555544e4c4c4d534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161616161616161616161616161616161616161616161616161616161616161616161615d554e4c4c4c535555554e4c4c4c534c4f555555514c4c55616161616161616161615b55514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555556606161616161616161615f4e51555555504c4c4c51576161616161616161616161554c4c51555555504c4c4c51555555504c4c4c5155555d61616161616161616161524c525555554f4c4c4c5257616161616161616161615d4c4c4c525555554f4c4c51616161616161616161615e554f4c4c4c525555554f4d5c616161616161616161616161616161616161616161616161616161616161616161616161616161616161615d554e4c4c4c535555554e4c4c4c534d4f545454514d4d55616161616161616161615b54514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545456606161616161616161615f4e50545454514d4d4d50566161616161616161616161554d4d50545454504d4d4d51545454504d4d4d5154545c61616161616161616161534d51545454504d4d4d5156616161616161616161615d4d4d4d51545454504d4d51616161616161616161615e54504d4d4d51545454504d5c616161616161616161616161616161616161616161616161616161616161616161616161616161616161615d544f4d4d4d525454544f4d4d4d5255514c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4f5f6161616161616161616056504c4c4c50555555504f60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616158554f4c4c4c515555554f50616161616161616161615e5555554f4c4c4c52555557616161616161616161615d4d525555554f4c4c4c52555e616161616161616161616161616161616161616161616161616161616161616161616161616161616161615a4c525555544e4c4c4c535555544e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e616161616161616161616161616161616161616161616161616161616161616161616161616161616161615a4c535555554e4c4c4c535555554e55524c4c4c5055555a61616161616161616161574c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4e5f6161616161616161616056504c4c4c51555555504e60616161616161616161615a5555504c4c4c51555555504c4c4c51555555504c4c596161616161616161616159554f4c4c4c525555554f4f616161616161616161615e5555554f4c4c4c52555558616161616161616161615d4d525555554f4c4c4c52555e616161616161616161616161616161616161616161616161616161616161616161616161616161616161615a4c535555554e4c4c4c535555554e54524d4d4d5054545a61616161616161616161584d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4f5f6161616161616161615f55514d4d4d50545454514f6061616161616161616161595454504d4d4d51545454504d4d4d51545454504d4d59616161616161616161615854504d4d4d515454545050616161616161616161615e545454504d4d4d51545457616161616161616161615d4d51545454504d4d4d51545e616161616161616161616161616161616161616161616161616161616161616161616161616161616161615a4d525454544f4d4d4d525454544f4c4f555555514c4c50585b5b5b59565656585b5855514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555658565656585b5b5b5956554d50555555504c4c4c50565b5b58565656595b5b5b58504c4c51555555504c4c4c51555555504c4c4c5155555958565656595b5b5b58564f4c515555554f4c4c4c52565b5b58565656595b5b5b564d4c4c525555554f4c4c4f595b5b5b57565656595b5a554f4c4c4c525555554f4d5356595b5b5b57565656595b5b5b57565656595b5b5b575656565a5b5b5b575656565a5b5b5b575656565a5b59544f4c4c4c535555544e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534d4f545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d515454544f4d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4d4d4d5255514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c515555554f4c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555544f4c4c4c525555544f4c4c4c525555544e4c4c4c535555544e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e54514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d50545454514d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4d4d4d525454544f4c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555544f4c4c4c525555544f4c4c4c535555544e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534d50545454514d4d3f2f313131302e2e2e2f313131302e2e2e2f313131302e2e2e2f313131302e2e2e30313131302e2e2e30313131302e2e2e30313131302e314c50545454514d4d4d505034312f2e2e2e303131312f414d4d51545454504d4d4d3d3131312f2e2e2e30313147504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d515454544a2e2e2e303131312f2e2e2e303131312f2e2e2e303131312f2e2e2e303131312f2f474d51545454504d4d4d513a31312f2e2e2e303131312f2e2e2e303131312f2e2e2e303131312f2e2e2e30313d544f4d4d4d525454544f4d4d4d5255514c4c4c5055553b1919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191f50504c4c4c5055555550461b191919191919191919193c5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c515555554f4c4c4c515555554f4c4c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2519191919191919191919191919191919191919191919191919191919191919192a4c525555544e4c4c4c535555544e55524c4c4c5055553b1919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191f51504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2419191919191919191919191919191919191919191919191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c5055553b1919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191f51504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2419191919191919191919191919191919191919191919191919191919191919192a4c535555554e4c4c4c535555554e54514d4d4d5054543b1919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191e4f514d4d4d5054545451471b191919191919191919193c5454504d4d4d515454542f191919191919191919193a51545454504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d451a191919191919191919191919191919191919191919191919191919191919191a4554504d4d4d51545454502519191919191919191919191919191919191919191919191919191919191919192a4d525454544f4d4d4d525454544f4c50555555514c4c361919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191e4851555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a191919191919191919191919191919191919191919191919191919191919191a404c525555554f4c4c4c522719191919191919191919191919191919191919191919191919191919191919192c554e4c4c4c535555554e4c4c4c534c4f555555514c4c361919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191e4851555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a191919191919191919191919191919191919191919191919191919191919191a3f4c525555554f4c4c4c522719191919191919191919191919191919191919191919191919191919191919192c554e4c4c4c535555554e4c4c4c534c4f555555514c4c361919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191e4851555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a191919191919191919191919191919191919191919191919191919191919191a3f4c525555554f4c4c4c522719191919191919191919191919191919191919191919191919191919191919192c554e4c4c4c535555554e4c4c4c534d4f545454514d4d371919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191e4a50545454514d4d4d504d1b19191919191919191919384d4d51545454504d4d4d2d191919191919191919193e504d4d4d51545454504d4d4d51545454504d4d4d51545454504d4d4d51545453461a191919191919191919191919191919191919191919191919191919191919191a414d51545454504d4d4d512619191919191919191919191919191919191919191919191919191919191919192c534f4d4d4d525454534f4d4d4d5255514c4c4c5055553b1919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191f50504c4c4c5155555550461b191919191919191919193c5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2519191919191919191919191919191919191919191919191919191919191919192a4c525555554e4c4c4c535555554e55524c4c4c5055553b1919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191919191f51504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2419191919191919191919191919191919191919191919191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c505555402121212121222222212121212122222221212121212119191919191919191919192121212122222221212121212222222121212121222751504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a1919191919191919191b2121212122222222212121212222222221212121222347554f4c4c4c525555554f2419191919191919191919212222222121212122222222212121212222222221212e4c535555554e4c4c4c535555554e54514d4d4d505454544f4c4c4c4e5151514f4c4c4c4e5151514f4c4c4c4e4c1c1919191919191919191b484c4c4e5151514e4c4c4c4e5151514e4c4c4c4e515153514d4d4d5054545451471b191919191919191919193b5454504d4d4d515454542f191919191919191919193a51545454504d4d4d51545454504d4d4d51545454504d4d4d51545453504d4d4d451a191919191919191919264e4c4c4c4f5151514e4c4c4c4f5151514e4c4c4c4f515254504d4d4d5154545450251919191919191919191b475151514d4c4c4c505151514d4c4c4c505151514d4c4c4d525454534f4d4d4d525454534f4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52271919191919191919191b434c4c4c525555554e4c4c4c525555554e4c4c4c525555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52271919191919191919191b434c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52271919191919191919191b434c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534e4f535353514e4e4e4f535353514e4e4e50535353514e4e4e5053535351491d1919191919191919191c4f5353514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504c1b19191919191919191919394e4e50535353504e4e4e2d191919191919191919193d504e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e50535353461a1919191919191919192451535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51261919191919191919191b444e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e525353534f4e4e4e5255514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193c5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f251919191919191919191a485555554e4c4c4c525555554e4c4c4c525555554e4c4c4c525555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f241919191919191919191a495555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f241919191919191919191a495555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e53524e4e4e4f535353514e4e4e4f535353514e4e4e50535353514e4e4e504e1e1919191919191919191b4a4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e5053535351481b191919191919191919193b5353504e4e4e515353532f191919191919191919193b51535353514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e451a19191919191919191925504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e5153535350251919191919191919191b47535353504e4e4e51535353504e4e4e51535353504e4e4e515353534f4e4e4e525353534f4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52271919191919191919191b434c4c4c525555554e4c4c4c525555554e4c4c4c525555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52271919191919191919191b434c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52271919191919191919191b434c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534e4f535353514e4e4e4f535353514e4e4e50535353514e4e4e5053535351491d1919191919191919191c4f5353514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504c1b19191919191919191919394e4e50535353504e4e4e2d191919191919191919193d504e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e50535353461a1919191919191919192451535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51261919191919191919191b444e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e525353534f4e4e4e5255514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c5155555550461b191919191919191919193c5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f251919191919191919191a485555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f241919191919191919191a495555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f241919191919191919191a495555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e53524e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504e1e1919191919191919191b4a4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e5053535351481b191919191919191919193b5353504e4e4e515353532f191919191919191919193b51535353514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e451a19191919191919191925504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e5153535350251919191919191919191b47535353504e4e4e51535353504e4e4e51535353504e4e4e515353534f4e4e4e515353534f4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c505555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52271919191919191919191b434c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52271919191919191919191b434c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52271919191919191919191b434c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534e4f535353514e4e4e50535353514e4e4e50535353514e4e4e5053535351491d1919191919191919191c4f5353514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504c1b19191919191919191919394e4e51535353504e4e4e2d191919191919191919193d504e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e50535353461a1919191919191919192451535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51261919191919191919191b444e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e515353534f4e4e4e5155514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c5155555550461b191919191919191919193c5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a1919191919191919192446434343484a4a4a46434343484a4a4a46434343484b54554f4c4c4c525555554f251919191919191919191a3f4a4a4a45434343484a4a4a45434343484a4a4a4543474c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2419191919191919191919191919191919191919191919191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2419191919191919191919191919191919191919191919191919191919191919192a4c535555554e4c4c4c535555554e53514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504d1e1919191919191919191b4a4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e5053535351481b191919191919191919193b5353504e4e4e515353532e191919191919191919193b51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e451a191919191919191919191919191919191919191919191919191919191919191a4453504e4e4e51535353502519191919191919191919191919191919191919191919191919191919191919192b4e515353534f4e4e4e525353534f4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c505555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a191919191919191919191919191919191919191919191919191919191919191a404c525555554f4c4c4c522719191919191919191919191919191919191919191919191919191919191919192c554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a191919191919191919191919191919191919191919191919191919191919191a3f4c525555554f4c4c4c522719191919191919191919191919191919191919191919191919191919191919192c554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a191919191919191919191919191919191919191919191919191919191919191a3f4c525555554f4c4c4c522719191919191919191919191919191919191919191919191919191919191919192c554e4c4c4c535555554e4c4c4c534e50535353514e4e4e50535353514e4e4e50535353514e4e4e5053535351491d1919191919191919191c4e5353514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504c1b19191919191919191919394e4e51535353504e4e4e2d191919191919191919193d504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353451a191919191919191919191919191919191919191919191919191919191919191a414e51535353504e4e4e512619191919191919191919191919191919191919191919191919191919191919192b534f4e4e4e525353534f4e4e4e5255514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c5155555550461b191919191919191919193c5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2519191919191919191919191919191919191919191919191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2419191919191919191919191919191919191919191919191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2419191919191919191919191919191919191919191919191919191919191919192a4c535555554e4c4c4c535555554e53514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504d1e1919191919191919191b4a4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e5053535351481b191919191919191919193b5353504e4e4e515353532e191919191919191919193b51535353504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e451a1919191919191919191b242525252423232324252525242323232425252524244653504e4e4e51535353502f2525242323232425252524232323242525252423231b191919191919191919192b4e515353534f4e4e4e525353534f4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924515353534d4b4b4b515353534d4b4b4b515353534d4b4c4c525555554f4c4c4c525453534d4b4b4b515353534d4b4b4b515353534d4b4b23191919191919191919192c554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c23191919191919191919192c554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c23191919191919191919192c554e4c4c4c535555554e4c4c4c534e50535353514e4e4e50535353514e4e4e50535353514e4e4e50535353514a1d1919191919191919191c4e5353504e4e4e50535353504e4e4e50535353514e4e4e50535353504e4e4e504c1b19191919191919191919394e4e51535353504e4e4e2d191919191919191919193d504e4e4e51535353504e4e4e51535353504e4e4e51535353504e4e4e51535352461a1919191919191919192451535352504e4e4e51535352504e4e4e51535353504e4e4e51535353504e4e4e515353534f4e4e4e515353534f4e4e4e51535353504e4e24191919191919191919192b52504e4e4e525353524f4e4e4e5255514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c53555525191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c53555525191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c53555525191919191919191919192a4c535555554e4c4c4c535555554e53514e4e4e50535353514e4e4e50535353514e4e4e50535353514e4e4e504d1e1919191919191919191b4b4e4e50535353504e4e4e50535353514e4e4e50535353504e4e4e5053535350481b191919191919191919193b5353504e4e4e515353532e191919191919191919193b51535353504e4e4e51535353504e4e4e51535353504e4e4e51535352504e4e4e451a19191919191919191925504e4e4e51535352504e4e4e51535352504e4e4e51535353504e4e4e51535353504e4e4e515353534f4e4e4e51535353504e4e4e51535325191919191919191919192b4e515353524f4e4e4e525353524f4c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c23191919191919191919192c554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c23191919191919191919192c554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c23191919191919191919192c554e4c4c4c535555554e4c4c4c534f4f525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514a1d1919191919191919191c4e5252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f504b1b19191919191919191919394f4f50525252514f4f4f2d191919191919191919193d504f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252461a1919191919191919192551525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f24191919191919191919192b52504f4f4f51525252504f4f4f5155514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c53555525191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c53555525191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c53555525191919191919191919192a4c535555554e4c4c4c535555554e52524f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f504d1e1919191919191919191b4b4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f5052525251481b191919191919191919193b5252504f4f4f505252522e191919191919191919193b50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f451a19191919191919191925504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525225191919191919191919192b4f51525252504f4f4f51525252504c50555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c505555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c23191919191919191919192c554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c23191919191919191919192c554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c191919191919191919193f504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c52555555451a19191919191919191924525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c23191919191919191919192c554e4c4c4c535555554e4c4c4c534f4f525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514a1d1919191919191919191c4e5252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f504b1b19191919191919191919394f4f50525252514f4f4f2d191919191919191919193d504f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252461a1919191919191919192551525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f24191919191919191919192b52504f4f4f51525252504f4f4f5155514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c53555525191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191939515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c461a191919191919191919264f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c53555525191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f19191919191919191919202728282827262626272828282726262627282828272d4c4c525555554f4c4c4c461a1919191919191919191c272626262728282827262626272828282726262627294c554f4c4c4c525555554f2f2626272828282626262627282828262626262728281b191919191919191919192a4c535555554e4c4c4c535555554e52524f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f504d1e1919191919191919191b4b4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f5052525251481b191919191919191919193a5252514f4f4f505252522e1919191919191919191919191919191919191919191919191919191919191919234f4f50525252514f4f4f451a191919191919191919191919191919191919191919191919191919191919191a4452504f4f4f51525252502519191919191919191919191919191919191919191919191919191919191919192b4f51525252504f4f4f51525252504c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c19191919191919191919191919191919191919191919191919191919191919192355554f4c4c4c52555555451a191919191919191919191919191919191919191919191919191919191919191a3f4c525555554f4c4c4c522719191919191919191919191919191919191919191919191919191919191919192c554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c19191919191919191919191919191919191919191919191919191919191919192355554f4c4c4c52555555451a191919191919191919191919191919191919191919191919191919191919191a3f4c525555554f4c4c4c522719191919191919191919191919191919191919191919191919191919191919192c554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551471d1919191919191919191c515555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c514e1b19191919191919191919374c4c51555555504c4c4c2c19191919191919191919191919191919191919191919191919191919191919192355554f4c4c4c52555555451a191919191919191919191919191919191919191919191919191919191919191a3f4c525555554f4c4c4c522719191919191919191919191919191919191919191919191919191919191919192c554e4c4c4c535555554e4c4c4c534f4f525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514a1d1919191919191919191c4e5252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f504b1b19191919191919191919394f4f50525252514f4f4f2d1919191919191919191919191919191919191919191919191919191919191919235252514f4f4f50525252461a191919191919191919191919191919191919191919191919191919191919191a424f51525252504f4f4f512619191919191919191919191919191919191919191919191919191919191919192b52504f4f4f51525252504f4f4f5155514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191919191919191919191919191919191919191919191919224c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2519191919191919191919191919191919191919191919191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191919191919191919191919191919191919191919191919224c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2419191919191919191919191919191919191919191919191919191919191919192a4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c504f1e1919191919191919191b484c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c5155555550461b191919191919191919193d5555504c4c4c515555552f1919191919191919191919191919191919191919191919191919191919191919224c4c525555554f4c4c4c461a191919191919191919191919191919191919191919191919191919191919191b46554f4c4c4c525555554f2419191919191919191919191919191919191919191919191919191919191919192a4c535555554e4c4c4c535555554e52514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f504d1e1919191919191919191b4b4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f5052525251491b191919191919191919193a5252504f4f4f515252522e1919191919191919191919191919191919191919191919191919191919191919234f4f50525252504f4f4f451a191919191919191919191919191919191919191919191919191919191919191a4352514f4f4f50525252512519191919191919191919191919191919191919191919191919191919191919192b4f51525252504f4f4f51525252504c4f555555514c4c4c50555555514c4c4c50555555514c4c4c5055555551481f1b1b1b1b1b1b1b1b1b1e515555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c514e1d1b1b1b1b1b1b1b1b1b1b384c4c51555555504c4c4c2e1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b2555554f4c4c4c52555555451c1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1c3f4c525555554f4c4c4c52281b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b1b2d554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4241444848484441414144535555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51544848444141414548484844474c4c51555555504c4c4c4948484844414141454848484441414145484848434141414548484843414141454955554f4c4c4c525555554f414141454848484341414146484848434141414648484843414141464848484341484c525555554f4c4c4c524a48484341414146484848434141414648484843414141464848484341414146484b554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f50525252514f4f4f50525252514f4f4f50525252504f4f4f50525252504f4f4f50525252504f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f5155524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e52514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252514f4f4f50525252514f4f4f50525252504f4f4f50525252504f4f4f50525252504f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534c4f555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c534f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f50525252514f4f4f50525252514f4f4f50525252514f4f4f50525251514f4f4f50525251514f4f4f50525251514f4f4f50525251514f4f4f50525252514f4f4f50525252514f4f4f50525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f51525252504f4f4f5155524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e55524c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555514c4c4c50555555504c4c4c50555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c51555555504c4c4c515555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c525555554f4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e4c4c4c535555554e;


always_ff @ (*) begin
	if ( DrawX >= start_x & DrawX < start_x + size_x & DrawY >= start_y & DrawY < start_y + size_y ) begin
		is_title <= 1'b1;
		data_R <= ROM_R[ (DrawY*234*2-:1) : (DrawY*234*2 + DrawX*2) ];
		DATA_OUT = char_font[2*ROW_NUM+:10]
		data_G <= ROM_G[ (DrawY*234*2 + DrawX*2 + 1) : (DrawY*234*2 + DrawX*2) ];
	end
	else begin
		is_title <= 1'b0;
		data_R <= 2'b00;
		data_G <= 2'b00;
	end
end
	
endmodule*/
