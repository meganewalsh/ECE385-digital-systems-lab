module testbench();

timeunit 10ns;	// Half clock cycle at 50 MHz
			// This is the amount of time represented by #1 
timeprecision 1ns;

// These signals are internal because the processor will be 
// instantiated as a submodule in testbench.
logic Clk = 0;
logic Reset, Run, ClearA_LoadB, X;
logic [7:0] S;
logic [7:0] Aval, Bval;
logic [6:0] AhexL, AhexU, BhexL, BhexU; 

// To store expected results
logic [7:0] ans_1a, ans_2b;
		
// Instantiating the DUT
// Make sure the module and signal names match with those in your design
top_level top_level0(.*);	

// Toggle the clock
// #1 means wait for a delay of 1 timeunit
always begin : CLOCK_GENERATION
#1 Clk = ~Clk;
end

initial begin: CLOCK_INITIALIZATION
    Clk = 0;
end 

// Testing begins here
// The initial block is not synthesizable
// Everything happens sequentially inside an initial block
// as in a software program
initial begin: TEST_VECTORS
Reset = 0;		// Toggle Rest
Reset = 1;
S = 8'b00000101;
ClearA_LoadB = 1;
S = 8'b00001111;
Run = 0;
Run = 1;
Run = 0;
Run = 1;
Run = 0;
Run = 1;
Run = 0;


end
endmodule
