module reg_x ();